`include "fourbyonemux.v"
module fourbyonemux_tb();
reg s0,s1,a1,b1,c1,d1;

wire out;

initial begin
$dumpfile("cmos_fourbyonemux.vcd");
$dumpvars(0,fourbyonemux_tb);
$display("s0,  s1,  in1,  in2,  in3,  in4,  out");
$monitor("%b,   %b,   %b,   %b,  %b,  %b,  %b", s0, s1, a1, b1, c1, d1, out);
#20 s0=0;s1=0;a1=0;b1=0;c1=0;d1=0;
#20 s0=0;s1=0;a1=0;b1=0;c1=0;d1=1;
#20 s0=0;s1=0;a1=0;b1=0;c1=1;d1=0;
#20 s0=0;s1=0;a1=0;b1=0;c1=1;d1=1;

#20 s0=0;s1=0;a1=0;b1=1;c1=0;d1=0;
#20 s0=0;s1=0;a1=0;b1=1;c1=0;d1=1;
#20 s0=0;s1=0;a1=0;b1=1;c1=1;d1=0;
#20 s0=0;s1=0;a1=0;b1=1;c1=1;d1=1;

#20 s0=0;s1=0;a1=1;b1=0;c1=0;d1=0;
#20 s0=0;s1=0;a1=1;b1=0;c1=0;d1=1;
#20 s0=0;s1=0;a1=1;b1=0;c1=1;d1=0;
#20 s0=0;s1=0;a1=1;b1=0;c1=1;d1=1;

#20 s0=0;s1=0;a1=1;b1=1;c1=0;d1=0;
#20 s0=0;s1=0;a1=1;b1=1;c1=0;d1=1;
#20 s0=0;s1=0;a1=1;b1=1;c1=1;d1=0;
#20 s0=0;s1=0;a1=1;b1=1;c1=1;d1=1;



#20 s0=0;s1=1;a1=0;b1=0;c1=0;d1=0;
#20 s0=0;s1=1;a1=0;b1=0;c1=0;d1=1;
#20 s0=0;s1=1;a1=0;b1=0;c1=1;d1=0;
#20 s0=0;s1=1;a1=0;b1=0;c1=1;d1=1;

#20 s0=0;s1=1;a1=0;b1=1;c1=0;d1=0;
#20 s0=0;s1=1;a1=0;b1=1;c1=0;d1=1;
#20 s0=0;s1=1;a1=0;b1=1;c1=1;d1=0;
#20 s0=0;s1=1;a1=0;b1=1;c1=1;d1=1;

#20 s0=0;s1=1;a1=1;b1=0;c1=0;d1=0;
#20 s0=0;s1=1;a1=1;b1=0;c1=0;d1=1;
#20 s0=0;s1=1;a1=1;b1=0;c1=1;d1=0;
#20 s0=0;s1=1;a1=1;b1=0;c1=1;d1=1;

#20 s0=0;s1=1;a1=1;b1=1;c1=0;d1=0;
#20 s0=0;s1=1;a1=1;b1=1;c1=0;d1=1;
#20 s0=0;s1=1;a1=1;b1=1;c1=1;d1=0;
#20 s0=0;s1=1;a1=1;b1=1;c1=1;d1=1;



#20 s0=1;s1=0;a1=0;b1=0;c1=0;d1=0;
#20 s0=1;s1=0;a1=0;b1=0;c1=0;d1=1;
#20 s0=1;s1=0;a1=0;b1=0;c1=1;d1=0;
#20 s0=1;s1=0;a1=0;b1=0;c1=1;d1=1;

#20 s0=1;s1=0;a1=0;b1=1;c1=0;d1=0;
#20 s0=1;s1=0;a1=0;b1=1;c1=0;d1=1;
#20 s0=1;s1=0;a1=0;b1=1;c1=1;d1=0;
#20 s0=1;s1=0;a1=0;b1=1;c1=1;d1=1;

#20 s0=1;s1=0;a1=1;b1=0;c1=0;d1=0;
#20 s0=1;s1=0;a1=1;b1=0;c1=0;d1=1;
#20 s0=1;s1=0;a1=1;b1=0;c1=1;d1=0;
#20 s0=1;s1=0;a1=1;b1=0;c1=1;d1=1;

#20 s0=1;s1=0;a1=1;b1=1;c1=0;d1=0;
#20 s0=1;s1=0;a1=1;b1=1;c1=0;d1=1;
#20 s0=1;s1=0;a1=1;b1=1;c1=1;d1=0;
#20 s0=1;s1=0;a1=1;b1=1;c1=1;d1=1;



#20 s0=1;s1=1;a1=0;b1=0;c1=0;d1=0;
#20 s0=1;s1=1;a1=0;b1=0;c1=0;d1=1;
#20 s0=1;s1=1;a1=0;b1=0;c1=1;d1=0;
#20 s0=1;s1=1;a1=0;b1=0;c1=1;d1=1;

#20 s0=1;s1=1;a1=0;b1=1;c1=0;d1=0;
#20 s0=1;s1=1;a1=0;b1=1;c1=0;d1=1;
#20 s0=1;s1=1;a1=0;b1=1;c1=1;d1=0;
#20 s0=1;s1=1;a1=0;b1=1;c1=1;d1=1;

#20 s0=1;s1=1;a1=1;b1=0;c1=0;d1=0;
#20 s0=1;s1=1;a1=1;b1=0;c1=0;d1=1;
#20 s0=1;s1=1;a1=1;b1=0;c1=1;d1=0;
#20 s0=1;s1=1;a1=1;b1=0;c1=1;d1=1;

#20 s0=1;s1=1;a1=1;b1=1;c1=0;d1=0;
#20 s0=1;s1=1;a1=1;b1=1;c1=0;d1=1;
#20 s0=1;s1=1;a1=1;b1=1;c1=1;d1=0;
#20 s0=1;s1=1;a1=1;b1=1;c1=1;d1=1;


#20 $finish;
end


cmos_fourbyonemux n(
.s0(s0),
.s1(s1),
.a(a1),
.b(b1),
.c(c1),
.d(d1),
.y(out)
);

endmodule
