$date
	Thu Aug 30 16:01:40 2018
$end
$version
	Icarus Verilog
$end
$timescale
	1s
$end
$scope module nortb $end
$var wire 1 ! out $end
$var reg 1 " a1 $end
$var reg 1 # b1 $end
$scope module n $end
$var wire 1 $ a $end
$var wire 1 % b $end
$var wire 1 & gnd $end
$var wire 1 ' vdd $end
$var wire 1 ( w $end
$var wire 1 ! y $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
x(
1'
0&
x%
x$
x#
x"
x!
$end
#20
0#
1!
1(
0%
0"
0$
#40
1"
0!
1$
#60
1#
z(
1%
0"
0!
0$
#80
1"
1$
#100
